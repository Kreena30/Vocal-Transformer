BZh91AY&SY�ȝ �_�Py���߰?���P~s���㮔A�DƦ� h �@ 4	"ja)梟�)��h�   ���zM�ODh     0&&�	�&L�&	���J�i)�4ɠ�jz��2�� 4�d�Q���A�\�0j���!V$�)"������@�tB�_��`�i m� TX��f+�)�&h���
jȄ���u�V����P#)���fM܊��6tOB��	�I�_�)�I"���uj�I��w����\`��5�9�A�55W����Pm��B�90=n���5��!X�ba�}�H��0�nc�ng<�#[���e:�6Wrc�	�$�}O`o�<bf���X�*3S�'(@S7O�$�,�QV��m��ѱ��D�[�'��`��".� 9��A
@r�e��e��gXB��^;�&"�T�|0Apا��`�~��z�C�3�`\��;B�*/JirБ	m�_~`5㈴��#�#8) ����>���>d�y!�G�y9_�����8���+-�)�֍�a5��v��c.��H��k�8h��P�#�i��B�DD1��e�
x@��ʘJU�n�0,%�Z>��B�)��t<�A1�,As�V�;d-L����8̑���
A�^������6%�#P���,:0CW�c��r3�D��JS6���+������.��)��K��Ӈ,��фh���2�������
��͉h	������P�Ɓ)W��@�.9
�v��knZ`b�4�I��k����U0(z��)['Y�k\ZbT���/lԇ`u�!��t�t=��5� ν�����(�hj�mݚU��a�$�bo��\t@;�7w�b�����c�;�1�b9���%t�(�[MRn��l����b��0D���;[VK�U���?NH[i1dS\.@�$��#����F��m��&�l�S�}��5�a �?nJ@�j�&~%p��ܑN$�r'@