BZh91AY&SY��w�  �_�Px���߰?���P>��p���QOj2�&Pf�j�Ѡ4z�ѓ���=M��  �   %4 �z(ڞSe=�zjm@ #F@0	����L&i��EjhS��T�MH�2a1\��H�
T�?w�W�46 �wy��œΚ�����,[�9vA��t�V�kV�h-a�2����)#�H ,ѹ�rDb#}Im�<�b��U� Ĕy��m�`�ٗT��Ab na�\�,��G%(Ca�EZ�K����GS�X�h����Ҕ�iBL��$��q��2�_Ւ�Y�H�y��	����,FN~��%��j(��e# �oa�9U�q���\��H���=t���0�~���E.�.�?�N���f�Jn���������r{��t�؜�A{Paf$FLYVԗX���v>��)5(�!`�&�B�rh�ݣ*y���0��]k�j�����ߒ4�KV�`}laFvU�{'��%dIŕ{H�4��a-F>�|E���hd���=D�x��{^��I�m�شҢ;���H�����_b��e_��kI��e�-jG������s5^5��s�n5�51��L�Ԣb3�,�d;lpW��I�43h�=���8��4fC\��\�ɇ��b"�v��� -�g�$�+�^[��&A��p�� ��j��ܭ��c+T˚���D�U�B�m��2Lߐ�a#0��pl���q��5��:�gLQ<bl$��*�֙ �+�1��,��OiT�"%��H����B��9D% lQtD3!�@H����@kX��]��BB�u�h